module pamPy #(
    parameter GENERAL_DATA_WIDTH = 8,
    parameter GENERAL_ADDR_WIDTH = 12,
    parameter GENERAL_ULA_WIDTH = 24,
    parameter GENERAL_INSTRUCTION_WIDTH = 16
    )(
        input general_clk, general_reset
    );

// block 1
wire [(GENERAL_ADDR_WIDTH-1):0] GENERAL_MUX_REG1_IN;                   // regJump
wire [(GENERAL_DATA_WIDTH-1):0] GENERAL_MUX_REG2_IN_0; // regArg
wire [(GENERAL_ADDR_WIDTH-1):0] GENERAL_MUX_REG2_IN_1; // tos
wire [(GENERAL_ADDR_WIDTH-1):0] GENERAL_MUX_REG2_IN_2; // pc
    // CONTROLS
wire [1:0] GENERAL_SEL_MUX_OP1, GENERAL_SEL_MUX_OP2;
wire GENERAL_CTRL_REG_OP1, GENERAL_CTRL_REG_OP2;
wire [3:0] GENERAL_SEL_ULA;
    //outputs
wire [(GENERAL_ULA_WIDTH-1):0] GENERAL_ULA_OUT;
wire GENERAL_REG_OVERFLOW_OUT, GENERAL_REG_COMP_OUT;
// ----------------------------------------------------------------------------
//block 2
wire [(GENERAL_ADDR_WIDTH-1):0] GENERAL_STACK_FUNCTION_OUT;
    // CONTROLS
wire GENERAL_CTRL_REG_ARG, GENERAL_CTRL_REG_INSTR, GENERAL_CTRL_REG_JUMP, GENERAL_CTRL_REG_PC, GENERAL_SEL_MUX_PC;
    //outputs
wire [(GENERAL_DATA_WIDTH-1):0] GENERAL_REG_ARG, GENERAL_REG_INSTR;
wire [(GENERAL_ADDR_WIDTH-1):0] GENERAL_REG_JUMP, GENERAL_REG_PC;
// ----------------------------------------------------------------------------
//block 3
wire [(GENERAL_ADDR_WIDTH-1):0] GENERAL_REG_TOS;
//controls
wire GENERAL_CTRL_REG_TOS_FUNCTION, GENERAL_SEL_SOMADOR_SUBTRATOR, GENERAL_CTRL_STACK_FUNCTION, GENERAL_CTRL_REG_DATA_RETURN;
//outputs
wire [(GENERAL_ADDR_WIDTH-1):0] GENERAL_STACK_TOS_OUT;
wire [(GENERAL_DATA_WIDTH-1):0] GENERAL_REG_DATA_RETURN_OUT;
// ----------------------------------------------------------------------------
// block 4
wire [(GENERAL_DATA_WIDTH-1):0] GENERAL_STACK_OUT;
//CONTROLS
wire [1:0] GENERAL_SEL_MUX_STACK, GENERAL_CTRL_REG_MEM_EXT, GENERAL_CTRL_REG_STACK;
wire GENERAL_SEL_MUX_TOS, GENERAL_CTRL_REG_TOS, GENERAL_CTRL_STACK, GENERAL_CTRL_MEM_EXT, GENERAL_CTRL_REG_ADDR;
// ----------------------------------------------------------------------------
BLOCK_ULA_OPS #(
    .DATA_WIDTH (GENERAL_DATA_WIDTH),
    .ADDR_WIDTH (GENERAL_ADDR_WIDTH),
    .ULA_WIDTH (GENERAL_ULA_WIDTH)
    ) block_1 (
        .clk (general_clk),
        .MUX_REG1_IN (GENERAL_MUX_REG1_IN),
        .REG1_IN (GENERAL_STACK_OUT_READ),
        .MUX_REG2_IN_0 (GENERAL_MUX_REG2_IN_0),
        .MUX_REG2_IN_1 (GENERAL_MUX_REG2_IN_1),
        .MUX_REG2_IN_2 (GENERAL_MUX_REG2_IN_2),
        .REG2_IN (GENERAL_STACK_OUT_READ),
        // CONTROLS
        .SEL_MUX1 (GENERAL_SEL_MUX_OP1),
        .SEL_MUX2 (GENERAL_SEL_MUX_OP2),
        .CTRL_REG_OP1 (GENERAL_CTRL_REG_OP1),
        .CTRL_REG_OP2 (GENERAL_CTRL_REG_OP2),
        .SEL_ULA (GENERAL_SEL_ULA),
        // OUTPUT
        .REG_COMP_OUT (GENERAL_REG_COMP_OUT),
        .REG_OVERFLOW_OUT (GENERAL_REG_OVERFLOW_OUT),
        .ULA_OUT (GENERAL_ULA_OUT)
        );

BLOCK_PC_INSTR_ARG #(
    .DATA_WIDTH (GENERAL_DATA_WIDTH),
    .ADDR_WIDTH (GENERAL_ADDR_WIDTH),
    .ULA_WIDTH (GENERAL_ULA_WIDTH),
    .INSTRUCTION_WIDTH (GENERAL_INSTRUCTION_WIDTH)
    ) block_2 (
            .clk (general_clk),
            .MUX_IN_0 (GENERAL_ULA_OUT),
            .MUX_IN_1 (GENERAL_STACK_FUNCTION_OUT),
            // CONTROLS
            .CTRL_REG_ARG (GENERAL_CTRL_REG_ARG),
            .CTRL_REG_INSTR (GENERAL_CTRL_REG_INSTR),
            .CTRL_REG_JUMP (GENERAL_CTRL_REG_JUMP),
            .CTRL_REG_PC (GENERAL_CTRL_REG_PC),
            .SEL_MUX (GENERAL_SEL_MUX_PC),
            //outputs
            .REG_ARG_OUT (GENERAL_REG_ARG),
            .REG_INSTR_OUT (GENERAL_REG_INSTR),
            .REG_JUMP_OUT (GENERAL_REG_JUMP),
            .REG_PC_OUT (GENERAL_REG_PC),
        );

BLOCK_FUNCTIONS #(
    .DATA_WIDTH (GENERAL_DATA_WIDTH),
    .ADDR_WIDTH (GENERAL_ADDR_WIDTH)
    ) block_3 (
        .clk (general_clk),
        .reset (general_reset),
        .STACK_FUNCTION_IN (GENERAL_REG_PC),
        .STACK_TOS_IN (GENERAL_REG_TOS),
        .REG_DATA_RETURN_IN (GENERAL_STACK_OUT),
        //CONTROLS
        .CTRL_REG_TOS_FUNCTION (GENERAL_CTRL_REG_TOS_FUNCTION),
        .CTRL_STACK_FUNCTION (GENERAL_CTRL_STACK_FUNCTION),
        .SEL_SOMADOR_SUBTRATOR (GENERAL_SEL_SOMADOR_SUBTRATOR),
        .CTRL_REG_DATA_RETURN (GENERAL_CTRL_REG_DATA_RETURN),
        //outputs
        .STACK_FUNCTION_OUT (GENERAL_STACK_FUNCTION_OUT),
        .STACK_TOS_OUT (GENERAL_STACK_TOS_OUT),
        .REG_DATA_RETURN_OUT (GENERAL_REG_DATA_RETURN_OUT)
    );

BLOCK_STACK_TOS #(
    .DATA_WIDTH (GENERAL_DATA_WIDTH),
    .ADDR_WIDTH (GENERAL_ADDR_WIDTH),
    .ULA_WIDTH (GENERAL_ULA_WIDTH)
    ) block_4 (
        .clk (general_clk),
        .reset (general_reset),
        .MUX_STACK_IN_0 (GENERAL_REG_ARG),
        .MUX_STACK_IN_2 (GENERAL_REG_DATA_RETURN_OUT),
        .MUX_STACK_TOS_IN_3 (GENERAL_ULA_OUT),
        .REG_ADDR_IN (GENERAL_REG_JUMP),
        .MUX_TOS_IN_1 (GENERAL_STACK_TOS_OUT),
        //controls
        .SEL_MUX_STACK (GENERAL_SEL_MUX_STACK),
        .SEL_MUX_TOS (GENERAL_SEL_MUX_TOS),
        .CTRL_REG_MEM_EXT (GENERAL_CTRL_REG_MEM_EXT),
        .CTRL_REG_STACK (GENERAL_CTRL_REG_STACK),
        .CTRL_REG_TOS (GENERAL_CTRL_REG_TOS),
        .CTRL_STACK (GENERAL_CTRL_STACK),
        .CTRL_MEM_EXT (GENERAL_CTRL_MEM_EXT),
        .CTRL_REG_ADDR (GENERAL_CTRL_REG_ADDR),
        //outputs
        .REG_STACK_OUT_READ (GENERAL_STACK_OUT_READ),
        .REG_TOS_OUT (GENERAL_MUX_REG2_IN_1)
    );
endmodule
